module button_controller (
	input i_clk,
	input i_button,
	output wire o_led
);

endmodule